library verilog;
use verilog.vl_types.all;
entity DV4_vlg_vec_tst is
end DV4_vlg_vec_tst;
